module ReadSlave();

endmodule
